module fa (
  input  logic input1,
  input  logic input2,
  input  logic carry_in,
  output logic sum,
  output logic carry_out
);

  // Your code here

endmodule
