module priority_encoder (
  input  logic [7:0] req,
  output logic [2:0] enc,
  output logic       valid
);

 // Your code here

endmodule
