module adder (
  input  logic [3:0] input1,
  input  logic [3:0] input2,
  input  logic       carry_in,
  output logic [3:0] sum,
  output logic       carry_out
);

  // Your code here


endmodule
